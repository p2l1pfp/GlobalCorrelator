library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity test_algo_array is
    port(
        clk1 : in STD_LOGIC;
        clk2 : in STD_LOGIC;
        data_in : in STD_LOGIC_VECTOR(31 downto 0);
        data_out : out STD_LOGIC_VECTOR(31 downto 0)
    );
end test_algo_array;

architecture Behavioral of test_algo_array is

    signal bram_to_hls : STD_LOGIC_VECTOR(63 downto 0);
    signal hls_to_ila : STD_LOGIC_VECTOR(31 downto 0);
    signal bram_address : STD_LOGIC_VECTOR(0 downto 0) := "0";
    
--    attribute mark_debug : string;
--    attribute mark_debug of bram_to_hls : signal is "true"; 

    component blk_mem_gen_0
    port(clka : IN STD_LOGIC;
        ena : IN STD_LOGIC;
        wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
        addra : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
        dina : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
        douta : OUT STD_LOGIC_VECTOR(63 DOWNTO 0));
    end component;

    component simple_algo_array_hw_0
    port(
        outA_V_Addr_A : OUT STD_LOGIC_VECTOR(31 downto 0);                
      --outA_V_address0 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0);     
        ap_start : IN STD_LOGIC;        
        ap_done : OUT STD_LOGIC;        
        ap_idle : OUT STD_LOGIC;        
        ap_ready : OUT STD_LOGIC;
        inA_V_Dout_A : IN STD_LOGIC_VECTOR(31 downto 0);       
        inB_V_Dout_A : IN STD_LOGIC_VECTOR(31 downto 0);
        outA_V_Din_A : out STD_LOGIC_VECTOR(31 downto 0));
       -- inA_V_q0 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
       -- inB_V_q0 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
       -- outA_V_d0 : OUT STD_LOGIC_VECTOR(31 DOWNTO 0));      
    end component;      

    component ila_0
    port(clk : IN STD_LOGIC;
        probe0 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        probe1 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        probe2 : IN STD_LOGIC_VECTOR(31 DOWNTO 0));
    end component;

begin

    --data_out <= x"00000000";

    process(clk1)
    begin
        if rising_edge(clk1) then
           
            --generate an address, just toggling between 1 and 0 
            -- (the current bram only has two addresses)
            if( bram_address = "1") then 
                bram_address <= "0"; 
            else
                bram_address <= "1";
            end if;
           
            data_out <= bram_to_hls(31 downto 0);

        end if; -- clk1 rising edge
    end process;

    
    my_bram_label : blk_mem_gen_0
        PORT MAP(
                clka  => clk1, 
                ena   => '1',
                wea   => "0", 
                addra => bram_address,
                dina  => x"0000000000000000", 
                douta => bram_to_hls);

    my_hls_label : simple_algo_array_hw_0
        PORT MAP(
                outA_V_Addr_A => open,  
                --outa_v_address0 => open,
                ap_start => '1',
                ap_done => open,
                ap_idle => open,
                ap_ready => open,
                inA_V_Dout_A => bram_to_hls(63 downto 32),
                inB_V_Dout_A => bram_to_hls(31 downto 0),
                outA_V_Din_A => hls_to_ila);
                --ina_v_q0 => bram_to_hls(63 downto 32),
                --inb_v_q0 => bram_to_hls(31 downto 0),
                --outa_v_d0 => hls_to_ila);
    
    my_ila_label : ila_0
        PORT MAP(
                clk => clk1,
                probe0 => bram_to_hls(63 downto 32),
                probe1 => bram_to_hls(31 downto 0),
                probe2 => hls_to_ila);
                    
    
end Behavioral;
